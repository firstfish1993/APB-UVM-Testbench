`include "uvm_macros.svh"
package coverage;
import uvm_pkg::*;
import rw_trans::*;

class apb_subscriber extends uvm_subscriber #(apb_rw);
    `uvm_component_utils(apb_subscriber)
  
    logic [31:0] addr;     //Address
    logic [31:0] data;     //Data - For write or read response
    logic apb_cmd;       //command type
    logic sel;
    logic enable; 
    logic ready;
  
    covergroup inputs;
      apb_addr: coverpoint addr {
	bins one_hot_bita[34] = {
	  32'h0000_0000,
	  32'h0000_0001,
	  32'h0000_0002,
	  32'h0000_0003,
	  32'h0000_0004,
	  32'h0000_0005,
	  32'h0000_0006,
	  32'h0000_0007,
	  32'h0000_0008,
	  32'h0000_0009,
	  32'h0000_000A,
	  32'h0000_000B,
	  32'h0000_000C,
	  32'h0000_000D,
	  32'h0000_000E,
	  32'h0000_000F
	}; 
      } 

      apb_data: coverpoint data {
	bins one_hot_bitb[34] = {
	  32'b0000_0000_0000_0000_0000_0000_0000_0000,
	  32'b0000_0000_0000_0000_0000_0000_0000_0001, 
	  32'b0000_0000_0000_0000_0000_0000_0000_0010, 
	  32'b0000_0000_0000_0000_0000_0000_0000_0100, 
	  32'b0000_0000_0000_0000_0000_0000_0000_1000, 
	  32'b0000_0000_0000_0000_0000_0000_0001_0000, 
	  32'b0000_0000_0000_0000_0000_0000_0010_0000, 
	  32'b0000_0000_0000_0000_0000_0000_0100_0000, 
	  32'b0000_0000_0000_0000_0000_0000_1000_0000, 
	  32'b0000_0000_0000_0000_0000_0001_0000_0000, 
	  32'b0000_0000_0000_0000_0000_0010_0000_0000, 
	  32'b0000_0000_0000_0000_0000_0100_0000_0000, 
	  32'b0000_0000_0000_0000_0000_1000_0000_0000, 
	  32'b0000_0000_0000_0000_0001_0000_0000_0000, 
	  32'b0000_0000_0000_0000_0010_0000_0000_0000, 
	  32'b0000_0000_0000_0000_0100_0000_0000_0000, 
	  32'b0000_0000_0000_0000_1000_0000_0000_0000, 
	  32'b0000_0000_0000_0001_0000_0000_0000_0000, 
	  32'b0000_0000_0000_0010_0000_0000_0000_0000, 
	  32'b0000_0000_0000_0100_0000_0000_0000_0000, 
	  32'b0000_0000_0000_1000_0000_0000_0000_0000, 
	  32'b0000_0000_0001_0000_0000_0000_0000_0000, 
	  32'b0000_0000_0010_0000_0000_0000_0000_0000, 
	  32'b0000_0000_0100_0000_0000_0000_0000_0000, 
	  32'b0000_0000_1000_0000_0000_0000_0000_0000, 
	  32'b0000_0001_0000_0000_0000_0000_0000_0000, 
	  32'b0000_0010_0000_0000_0000_0000_0000_0000, 
	  32'b0000_0100_0000_0000_0000_0000_0000_0000, 
	  32'b0000_1000_0000_0000_0000_0000_0000_0000, 
	  32'b0001_0000_0000_0000_0000_0000_0000_0000, 
	  32'b0010_0000_0000_0000_0000_0000_0000_0000, 
	  32'b0100_0000_0000_0000_0000_0000_0000_0000, 
	  32'b1000_0000_0000_0000_0000_0000_0000_0000,  
	  32'b1111_1111_1111_1111_1111_1111_1111_1111 
	}; 
      }

      apb_cross: cross apb_addr, apb_data, apb_cmd;    
    endgroup
    
  function new(string name, uvm_component parent);
    super.new(name,parent);
    inputs=new;
  endfunction: new

  function void write(apb_rw t);
    addr = {t.addr};
    data = {t.data};
    apb_cmd = {t.apb_cmd};
    sel = {t.sel};
    enable = {t.enable};
    ready = {t.ready};
    inputs.sample();
  endfunction: write
endclass

endpackage: coverage
